module attack