module config

pub const (
	//Colors
    default          = "\x1b[39m"
    black            = "\x1b[30m"
    red              = "\x1b[31m"
    green            = "\x1b[32m"
    yellow           = "\x1b[33m"
    blue             = "\x1b[34m"
    purple           = "\x1b[35m"
    cyan             = "\x1b[36m"
    light_grey       = "\x1b[37m"
    dark_grey        = "\x1b[90m"
    light_red        = "\x1b[91m"
    light_green      = "\x1b[92m"
    light_yellow     = "\x1b[93m"
    light_blue       = "\x1b[94m"
    light_purple     = "\x1b[95m"
    light_cyan       = "\x1b[96m"
    white            = "\x1b[97m"
    // Background Colors
    default_bg       = "\x1b[49m"
    black_bg         = "\x1b[40m"
    red_bg           = "\x1b[41m"
    green_bg         = "\x1b[42m"
    yellow_bg        = "\x1b[43m"
    blue_bg          = "\x1b[44m"
    purple_bg        = "\x1b[45m"
    cyan_bg          = "\x1b[46m"
    light_gray_bg    = "\x1b[47m"
    dark_gray_bg     = "\x1b[100m"
    light_red_bg     = "\x1b[101m"
    light_green_bg   = "\x1b[102m"
    light_yellow_bg  = "\x1b[103m"
    light_blue_bg    = "\x1b[104m"
    light_purple_bg  = "\x1b[105m"
    light_cyan_bg    = "\x1b[106m"
    white_bg         = "\x1b[107m"
	// Extra ANSI Shit
	clear			 = "\033[2J\033[1;1H"
)