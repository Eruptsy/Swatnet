module logger