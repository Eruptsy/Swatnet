module api

import vweb
