module attack

pub fn send_api_attack(mut a AttackInfo) {
	
}