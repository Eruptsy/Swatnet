module cnc