module auth


// pub fn user_auth(usern string, passw string) string {
// 	mut c := crud.User{}
// }